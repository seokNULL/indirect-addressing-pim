module aim_subsys_top_wrapper #
  (
      parameter integer AXI_ID_WIDTH     = 2,
      parameter integer AXI_MASK_WIDTH   = 16,
      parameter integer AXI_DATA_WIDTH   = 256,
      parameter integer AXI_ADDR_WIDTH   = 32,
      parameter integer AXI_AWUSER_WIDTH = 0,
      parameter integer AXI_ARUSER_WIDTH = 0,
      parameter integer AXI_WUSER_WIDTH  = 0,
      parameter integer AXI_RUSER_WIDTH  = 0,
      parameter integer AXI_BUSER_WIDTH  = 0,
      parameter integer ADDR_LSB         = $clog2(AXI_DATA_WIDTH) - 3,
      parameter integer RD_DATA_DEPTH    = 64,
      parameter integer CH_NUM           = 3
  )
  (
  input                          sys_clk_n,
  input                          sys_clk_p,
  input                          sys_rst,
  output                         aclk,
  output                         clk_mcs,
  output                         rst_mcs,
  // AXI4: Write Address Channel
  input   [AXI_ID_WIDTH-1:0]     s_axi_awid,
  input   [AXI_ADDR_WIDTH-1:0]   s_axi_awaddr,
  input   [7:0]                  s_axi_awlen,
  input   [2:0]                  s_axi_awsize,
  input   [1:0]                  s_axi_awburst,
  input                          s_axi_awlock,
  input   [3:0]                  s_axi_awcache,
  input   [2:0]                  s_axi_awprot,
  input   [3:0]                  s_axi_awqos,
  input   [3:0]                  s_axi_awregion,
  input                          s_axi_awvalid,
  output                         s_axi_awready,
  // AXI4: Write Data Channel
  input   [AXI_DATA_WIDTH-1:0]   s_axi_wdata,
  input   [AXI_DATA_WIDTH/8-1:0] s_axi_wstrb,
  input                          s_axi_wlast,
  input                          s_axi_wvalid,
  output                         s_axi_wready,
  // AXI4: Write Response Channel
  output  [AXI_ID_WIDTH-1:0]     s_axi_bid,
  output  [1:0]                  s_axi_bresp,
  output                         s_axi_bvalid,
  input                          s_axi_bready,
  // AXI4: Read Address Channel
  input   [AXI_ID_WIDTH-1:0]     s_axi_arid,
  input   [AXI_ADDR_WIDTH-1:0]   s_axi_araddr,
  input   [7:0]                  s_axi_arlen,
  input   [2:0]                  s_axi_arsize,
  input   [1:0]                  s_axi_arburst,
  input                          s_axi_arlock,
  input   [3:0]                  s_axi_arcache,
  input   [2:0]                  s_axi_arprot,
  input   [3:0]                  s_axi_arqos,
  input   [3:0]                  s_axi_arregion,
  input                          s_axi_arvalid,
  output                         s_axi_arready,
  // AXI4: Read Data Channel
  output  [AXI_ID_WIDTH-1:0]     s_axi_rid,
  output  [AXI_DATA_WIDTH-1:0]   s_axi_rdata,
  output  [1:0]                  s_axi_rresp,
  output                         s_axi_rlast,
  output                         s_axi_rvalid,
  input                          s_axi_rready,
  // MCS IO Interface
  input                          IO_addr_strobe,
  input                          IO_read_strobe,
  input                          IO_write_strobe,
  input   [31:0]                 IO_address,
  input   [3:0]                  IO_byte_enable,
  input   [31:0]                 IO_write_data,
  output  [31:0]                 IO_read_data,
  output                         IO_ready,
  // LED Interface
  output  [CH_NUM-1:0]           led,

  // AiM (GDDR6) Interface
  output  [((CH_NUM-1)>>1):0]    CK_t, 
  output  [((CH_NUM-1)>>1):0]    CK_c,
  output  [((CH_NUM-1)>>1):0]    RESET_n,
  output  [CH_NUM-1:0] [9:0]     CA,
  output  [CH_NUM-1:0]           CABI_n,
  output  [CH_NUM-1:0]           CKE_n,
  output  [CH_NUM-1:0]           WCK1_t,
  output  [CH_NUM-1:0]           WCK1_c,
  output  [CH_NUM-1:0]           WCK0_t,
  output  [CH_NUM-1:0]           WCK0_c,
  inout  tri   [CH_NUM-1:0] [15:0]    DQ,

  inout  tri   [CH_NUM-1:0] [1:0]     EDC
  );


aim_subsys U0_AIM_SUBSYS(

 .sys_clk_n (sys_clk_n),
 .sys_clk_p (sys_clk_p),
 .sys_rst (sys_rst),
 .aclk (aclk),
 .clk_mcs (clk_mcs),
 .rst_mcs (rst_mcs),
 // AXI4: Write Address Channel
 .s_axi_awid (s_axi_awid),
 .s_axi_awaddr (s_axi_awaddr),
 .s_axi_awlen (s_axi_awlen),
 .s_axi_awsize (s_axi_awsize),
 .s_axi_awburst (s_axi_awburst),
 .s_axi_awlock (s_axi_awlock),
 .s_axi_awcache (s_axi_awcache),
 .s_axi_awprot (s_axi_awprot),
 .s_axi_awqos (s_axi_awqos),
 .s_axi_awregion (s_axi_awregion),
 .s_axi_awvalid (s_axi_awvalid),
 .s_axi_awready (s_axi_awready),
 // AXI4: Write Data Channel
 .s_axi_wdata (s_axi_wdata),
 .s_axi_wstrb (s_axi_wstrb),
 .s_axi_wlast (s_axi_wlast),
 .s_axi_wvalid (s_axi_wvalid),
 .s_axi_wready (s_axi_wready),
 // AXI4: Write Response Channel
 .s_axi_bid (s_axi_bid),
 .s_axi_bresp (s_axi_bresp),
 .s_axi_bvalid (s_axi_bvalid),
 .s_axi_bready (s_axi_bready),
 // AXI4: Read Address Channel
 .s_axi_arid (s_axi_arid),
 .s_axi_araddr (s_axi_araddr),
 .s_axi_arlen (s_axi_arlen),
 .s_axi_arsize (s_axi_arsize),
 .s_axi_arburst (s_axi_arburst),
 .s_axi_arlock (s_axi_arlock),
 .s_axi_arcache (s_axi_arcache),
 .s_axi_arprot (s_axi_arprot),
 .s_axi_arqos (s_axi_arqos),
 .s_axi_arregion (s_axi_arregion),
 .s_axi_arvalid (s_axi_arvalid),
 .s_axi_arready (s_axi_arready),
 // AXI4: Read Data Channel
 .s_axi_rid (s_axi_rid),
 .s_axi_rdata (s_axi_rdata),
 .s_axi_rresp (s_axi_rresp),
 .s_axi_rlast (s_axi_rlast),
 .s_axi_rvalid (s_axi_rvalid),
 .s_axi_rready (s_axi_rready),
 // MCS IO Interface
 .IO_addr_strobe (IO_addr_strobe),
 .IO_read_strobe (IO_read_strobe),
 .IO_write_strobe (IO_write_strobe),
 .IO_address (IO_address),
 .IO_byte_enable (IO_byte_enable),
 .IO_write_data (IO_write_data),
 .IO_read_data (IO_read_data),
 .IO_ready (IO_ready),
 // LED Interface
 .led (led),
 // AiM (GDDR6) Interface
 .CK_t (CK_t),
 .CK_c (CK_c),
 .RESET_n (RESET_n),
 .CA (CA),
 .CABI_n (CABI_n),
 .CKE_n (CKE_n),
 .WCK1_t (WCK1_t),
 .WCK1_c (WCK1_c),
 .WCK0_t (WCK0_t),
 .WCK0_c (WCK0_c),
 .DQ (DQ),
 .EDC (EDC)

);

endmodule